module tb_initial_message;

    initial begin
        $display("System Initialization Started...");
    end
endmodule