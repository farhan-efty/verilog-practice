int temperatures [] = '{-32, 45, 28, 50, 41, 39, 30};
int below_freezing [] = temperatures.find(x) with (x<0);

$display("Temperatures below freezing: %p", below_freezing);
