typedef struct packed {
    logic    RX_FLUSH;
    logic    TX_FLUSH;
    logic    CLK_EN;
} ctrl_reg_t;